// Code your testbench here
// or browse Examples
`include "uvm_pkg.sv"
import uvm_pkg::*;



`include "axi_global_usage.sv"
`include "interface.sv"

`include "axi_seq_item.sv"
`include "axi_seq.sv"
`include "axi_sqr.sv"
`include "axi_drv.sv"
`include "axi_mon.sv"
`include "axi_resp.sv"
`include "axi_agent.sv"
`include "axi_sco.sv"
`include "axi_cov.sv"

`include "axi_env.sv"
`include "axi_test.sv"
`include "testbench_top.sv"
