class axi_sqr extends uvm_sequencer#(axi_seq_item);
	`uvm_component_utils(axi_sqr)

  `UVM_COMP

endclass
